module microcode(
    input [15:0] reg_out,
	output reg [1:0] condition,
	output reg BT,
	output reg [48:0] OPs,
	output reg [6:0] jump_addr
); 
	
reg [58:0] ucode [0:75];
		
initial 
    begin
		ucode[0] = {3'b000,7'd1,49'd274877906944};
		ucode[1] = {3'b000,7'd2,49'd67108866};
		ucode[2] = {3'b100,7'd0,49'd141012366262272};
		ucode[3] = {3'b000,7'd4,49'd67108866};
		ucode[4] = {3'b000,7'd5,49'd549755813888};
		ucode[5] = {3'b000,7'd6,49'd1};
		ucode[6] = {3'b000,7'd0,49'd128};
		ucode[7] = {3'b000,7'd8,49'd67108866};
		ucode[8] = {3'b000,7'd9,49'd549755813888};
		ucode[9] = {3'b000,7'd10,49'd1};
		ucode[10] = {3'b000,7'd0,49'd16};
		ucode[11] = {3'b000,7'd12,49'd137438953472};
		ucode[12] = {3'b000,7'd13,49'd131072};
		ucode[13] = {3'b000,7'd14,49'd512};
		ucode[14] = {3'b000,7'd0,49'd2048};
		ucode[15] = {3'b000,7'd16,49'd137438953472};
		ucode[16] = {3'b000,7'd17,49'd2097152};
		ucode[17] = {3'b000,7'd18,49'd512};
		ucode[18] = {3'b000,7'd19,49'd4294967296};
		ucode[19] = {3'b000,7'd0,49'd16777216};
		ucode[20] = {3'b000,7'd21,49'd137438953472};
		ucode[21] = {3'b000,7'd22,49'd131072};
		ucode[22] = {3'b000,7'd23,49'd512};
		ucode[23] = {3'b000,7'd24,49'd2097152};
		ucode[24] = {3'b000,7'd25,49'd17179869184};
		ucode[25] = {3'b000,7'd26,49'd4294967296};
		ucode[26] = {3'b000,7'd27,49'd4294967296};
		ucode[27] = {3'b000,7'd0,49'd16448};
		ucode[28] = {3'b000,7'd29,49'd137438953472};
		ucode[29] = {3'b000,7'd30,49'd262144};
		ucode[30] = {3'b000,7'd31,49'd17592186044416};
		ucode[31] = {3'b000,7'd32,49'd8192};
		ucode[32] = {3'b000,7'd33,49'd137438953472};
		ucode[33] = {3'b000,7'd34,49'd35184372088832};
		ucode[34] = {3'b000,7'd35,49'd1048576};
		ucode[35] = {3'b000,7'd36,49'd17179869184};
		ucode[36] = {3'b000,7'd0,49'd281474976776192};
		ucode[37] = {3'b000,7'd38,49'd524288};
		ucode[38] = {3'b000,7'd39,49'd8589934592};
		ucode[39] = {3'b000,7'd40,49'd512};
		ucode[40] = {3'b000,7'd0,49'd2199023255552};
		ucode[41] = {3'b000,7'd42,49'd8589934592};
		ucode[42] = {3'b000,7'd43,49'd2148007936};
		ucode[43] = {3'b000,7'd44,49'd512};
		ucode[44] = {3'b000,7'd0,49'd8796093022208};
		ucode[45] = {3'b000,7'd46,49'd1073741856};
		ucode[46] = {3'b000,7'd47,49'd1};
		ucode[47] = {3'b000,7'd0,49'd134217728};
		ucode[48] = {3'b000,7'd49,49'd536870912};
		ucode[49] = {3'b000,7'd50,49'd1};
		ucode[50] = {3'b000,7'd0,49'd134217728};
		ucode[51] = {3'b000,7'd52,49'd268435456};
		ucode[52] = {3'b000,7'd53,49'd1};
		ucode[53] = {3'b000,7'd0,49'd134217728};
		ucode[54] = {3'b000,7'd0,49'd137438953472};
		ucode[55] = {3'b000,7'd0,49'd34359738368};
		ucode[56] = {3'b000,7'd0,49'd4194304};
		ucode[57] = {3'b000,7'd0,49'd8192};
		ucode[58] = {3'b000,7'd0,49'd8425472};
		ucode[59] = {3'b000,7'd0,49'd2097152};
		ucode[60] = {3'b000,7'd0,49'd131072};
		ucode[61] = {3'b000,7'd0,49'd4466765987840};
		ucode[62] = {3'b000,7'd0,49'd1048576};
		ucode[63] = {3'b000,7'd64,49'd268500992};
		ucode[64] = {3'b000,7'd65,49'd4};
		ucode[65] = {3'b000,7'd0,49'd1280};
		ucode[66] = {3'b001,7'd69,49'd0};
		ucode[67] = {3'b000,7'd68,49'd2};
		ucode[68] = {3'b000,7'd0,49'd33554432};
		ucode[69] = {3'b000,7'd0,49'd67108864};
		ucode[70] = {3'b000,7'd0,49'd70368744177664};
		ucode[71] = {3'b000,7'd0,49'd1099511627776};
		ucode[72] = {3'b000,7'd0,49'd512};
		ucode[73] = {3'b000,7'd0,49'd17179869184};
		ucode[74] = {3'b000,7'd0,49'd8};
		ucode[75] = {3'b000,7'd0,49'd35184372088840}; // new line

	end

//Issuing first micro code at the start
initial {BT, condition, jump_addr, OPs} = ucode[0];
	
always @(reg_out)
	{BT, condition, jump_addr, OPs}= ucode[reg_out];
			
endmodule